library ieee;
    use ieee.std_logic_1164.all;

package p_axi is

  type axi_s_d1 is record
     tdata  : std_logic_vector(8 -1 downto 0);
     tlast  : std_logic;
     tvalid : std_logic; 
     tuser  : std_logic;
  end record;

  type axi_s_d2 is record
     tready : std_logic;
  end record;

end package;

package body p_axi is

end p_axi;